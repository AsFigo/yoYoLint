/*
module two_2d_arr #(
     parameter WDT = 3,
     parameter CNT = 2
) (
     input [WDT-1:0] in_a [CNT-1:0],
     output [WDT-1:0] out_b [CNT-1:0]
);
endmodule
*/
module top(output int a, b, c, d);
/*
   int x [3:0] = '{10, 11, 12, 13};

   assign a = x[0];
   assign b = x[1];
   assign c = x[2];
   assign d = x[3];
   */
endmodule

