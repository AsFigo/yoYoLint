package my_pkg;
      parameter KL=64;
endpackage


import my_pkg::*;
module top(
    input logic i_clk,
    output logic o_done
);
endmodule